module test(input logic A, clk, output logic B);
	assign A = B;
endmodule
